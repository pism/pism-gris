netcdf pism_overrides {
    variables:
    byte pism_overrides;

    pism_overrides:stress_balance.sia.max_diffusivity = 100000.0;
    pism_overrides:stress_balance.sia.max_diffusivity_doc = "Maximum allowed diffusivity of the SIA flow. PISM stops with an error message if the SIA diffusivity exceeds this limit.";
    pism_overrides:stress_balance.sia.max_diffusivity_type = "scalar";
    pism_overrides:stress_balance.sia.max_diffusivity_units = "m2 s-1";

    pism_overrides:surface.pdd.air_temp_all_precip_as_snow = 272.15;
    pism_overrides:surface.pdd.air_temp_all_precip_as_snow_doc = "Kelvin; threshold temperature below which all precipitation is snow";

    pism_overrides:surface.pdd.air_temp_all_precip_as_rain = 274.15;
    pism_overrides:surface.pdd.air_temp_all_precip_as_rain_doc = "Kelvin; threshold temperature above which all precipitation is rain; must exceed air_temp_all_precip_as_snow to avoid division by zero, because difference is in a denominator";

    pism_overrides:surface.pdd.refreeze = 0.47;
    pism_overrides:surface.pdd.refreeze_doc = "EISMINT-Greenland value [@ref RitzEISMINT]";
    pism_overrides:surface.pdd.refreeze_type = "scalar";
    pism_overrides:surface.pdd.refreeze_units = "1";

    pism_overrides:surface.pdd.refreeze_ice_melt = "no";
    pism_overrides:surface.pdd.refreeze_ice_melt_doc = "If set to 'yes', refreeze surface.pdd.refreeze fraction of melted ice, otherwise all of the melted ice runs off.";
    pism_overrides:surface.pdd.refreeze_ice_melt_type = "boolean";

    pism_overrides:run_info.institution = "University of Alaska Fairbanks";
    pism_overrides:run_info.institution_doc = "Institution name. This string is written to output files as the 'institution' global attribute.";

    pism_overrides:output.backup_interval = 5.0;
    pism_overrides:output.backup_interval_doc = "hours; wall-clock time between automatic backups";
    
    pism_overrides:surface.force_to_thickness.alpha = 1.0;
    pism_overrides:surface.force_to_thickness.alpha_doc = "yr-1; exponential coefficient in force-to-thickness mechanism";

    pism_overrides:surface.force_to_thickness.ice_free_alpha_factor = 10.0;
    pism_overrides:surface.force_to_thickness.ice_free_alpha_factor_doc = "; force_to_thickness_alpha is multiplied by this factor in areas that are ice-free according to the target ice thickness and force_to_thickness_ice_free_thickness_threshold";

    pism_overrides:ocean.sub_shelf_heat_flux_into_ice = 50.0;
    pism_overrides:ocean.sub_shelf_heat_flux_into_ice_doc = "W m-2; = J m-2 s-1; naively chosen default value for heat from ocean; see comments in @ref pism::POConstant::shelf_base_mass_flux().";

    pism_overrides:climate_forcing.buffer_size = 13;
    pism_overrides:climate_forcing.buffer_size_doc = "; number of 2D climate forcing records to keep in memory; = 5 years of monthly records";

    pism_overrides:geometry.ice_free_thickness_standard_units = "meters";
    pism_overrides:geometry.ice_free_thickness_standard_type = "scalar";
    pism_overrides:geometry.ice_free_thickness_standard = 10.0;
    pism_overrides:geometry.ice_free_thickness_standard_doc = "If ice is thinner than this standard then the mask is set to MASK_ICE_FREE_BEDROCK or MASK_ICE_FREE_OCEAN.";

}
